module mem_cycle();




always @(posedge clock)
begin


end

endmodule