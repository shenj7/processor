// module forward_unit_component();

// input clock;
// input memread;

// output reg write;

// always @(posedge clock)
// begin
//     //0 if we want to stall otherwise 1 (should mostly be 1)
//     if (memread == 1) begin
//         stall = 0;
//     end else begin
//         stall = 1;
//     end
// end



// endmodule