module load_store(clock, read_in, rst, write_out);

endmodule