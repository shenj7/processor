//replace inst mem in load_store.v

module inst_mem_wrapper();




endmodule